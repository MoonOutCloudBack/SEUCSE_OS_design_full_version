// 用来显示 shell 的 vga 模块
// 魔改了 https://www.cnblogs.com/liujinggang/p/9690504.html 的框架


module mfp_ahb_vga_shell_output(
    input                   I_clk   ,       // 系统 50MHz 时钟
    input                   I_rst_n ,       // 系统复位
    
    input           [12287:0]  I_string,    // 希望显示的字符串，64 * 24 * 8 = 12288
    output  reg     [3:0]    O_red   ,      // VGA 红色分量
    output  reg     [3:0]    O_green ,      // VGA 绿色分量
    output  reg     [3:0]    O_blue  ,      // VGA 蓝色分量
    output                  O_hs    ,       // VGA 行同步信号
    output                  O_vs            // VGA 场同步信号
    // 共 14 个输出信号
);
    
    
    // 关于 VGA 的时序信号：
    // 可参考 https://blog.csdn.net/u014586651/article/details/121850814
    // 行时序：
        // 包括：行同步 (Hor Sync)、行消隐 (Hor Back Porch)、行视频有效 (Hor Active Video)、行前肩 (Hor Front Porch)
        // 在一个行周期内，行时序输出首先在 行同步 时间内置零，然后保持 1。
        // 数据输出：首先等一个 行消隐，然后在 行视频有效 时间段内输出，最后等一个 行前肩
    // 场时序：
        // 包括：场同步 (Ver Sync)、场消隐 (Ver Back Porch)、场视频有效 (Ver Active Video)、场前肩 (Ver Front Porch)
        // 在一个场周期内，场时序输出首先在 场同步 时间内置零，然后保持 1。
        // 数据输出：首先等一个 场消隐，然后在 场视频有效 时间段内输出，最后等一个 场前肩
    // 需要注意：
        // 行时序以 像素 为单位， 场时序以 行 为单位
        // 分辨率为 640*480 时，要用 25.275 MHz 的时钟

    
    // 关于 VGA 同步 shell 输出：
        // 字模：
            // 一行有 640 个像素，要摆 64 个字符，一个字符 10 像素
            // 一列有 480 个像素，要摆 24 个字符，一个字符 20 像素
            // 因此，使用比例为 1：2 的字模
        // 判断当前为哪个字符：
            // 用行计数器得到 x 坐标，场计数器得到 y 坐标，直接索引输入字符串
        // 输出字模：
            // 只找到了 8 * 16 的字模，因此边缘留白
            // 用像素在 10 * 20 字符里的 x y 坐标，索引字模 parameter

    
    // 分辨率为 640*480 时，行时序各个参数定义
    parameter       C_H_SYNC_PULSE      =   96  , 
                    C_H_BACK_PORCH      =   48  ,
                    C_H_ACTIVE_TIME     =   640 ,
                    C_H_FRONT_PORCH     =   16  ,
                    C_H_LINE_PERIOD     =   800 ;

    // 分辨率为 640*480 时，场时序各个参数定义               
    parameter       C_V_SYNC_PULSE      =   2   , 
                    C_V_BACK_PORCH      =   33  ,
                    C_V_ACTIVE_TIME     =   480 ,
                    C_V_FRONT_PORCH     =   10  ,
                    C_V_FRAME_PERIOD    =   525 ;
                    
    reg [11:0]      R_h_cnt         ; // 行时序计数器
    reg [11:0]      R_v_cnt         ; // 列时序计数器
    reg             R_clk_25M       ; // 25MHz 像素时钟

    wire            W_active_flag   ; // 激活标志，当这个信号为 1 时 RGB 的数据可以显示在屏幕上

    // 为了输出 shell 的自定义 reg 变量
    reg [5:0]       R_char_h_cnt    ; // 打印字符的当前行坐标
    reg [4:0]       R_char_v_cnt    ; // 打印字符的当前列坐标
    reg [7:0]       R_now_ascii     ; // 打印字符的 8 位 ASCII 码
    reg [3:0]       R_char_h_detail ; // 打印字符 字模的当前行坐标
    reg [4:0]       R_char_v_detail ; // 打印字符 字模的当前列坐标

    // 133 * 16 * 8 字模的 parameter
    parameter [7:0] C_ascii_character [2127:0] =
    {   
        0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,       //0x00
        0x00,0x00,0x7E,0x81,0xA5,0x81,0x81,0xBD,0x99,0x81,0x81,0x7E,0x00,0x00,0x00,0x00,       //0x01
        0x00,0x00,0x7E,0xFF,0xDB,0xFF,0xFF,0xC3,0xE7,0xFF,0xFF,0x7E,0x00,0x00,0x00,0x00,       //0x02
        0x00,0x00,0x00,0x00,0x6C,0xFE,0xFE,0xFE,0xFE,0x7C,0x38,0x10,0x00,0x00,0x00,0x00,       //0x03
        0x00,0x00,0x00,0x00,0x10,0x38,0x7C,0xFE,0x7C,0x38,0x10,0x00,0x00,0x00,0x00,0x00,       //0x04
        0x00,0x00,0x00,0x18,0x3C,0x3C,0xE7,0xE7,0xE7,0x18,0x18,0x3C,0x00,0x00,0x00,0x00,       //0x05
        0x00,0x00,0x00,0x18,0x3C,0x7E,0xFF,0xFF,0x7E,0x18,0x18,0x3C,0x00,0x00,0x00,0x00,       //0x06
        0x00,0x00,0x00,0x00,0x00,0x00,0x18,0x3C,0x3C,0x18,0x00,0x00,0x00,0x00,0x00,0x00,       //0x07
        0xFF,0xFF,0xFF,0xFF,0xFF,0xFF,0xE7,0xC3,0xC3,0xE7,0xFF,0xFF,0xFF,0xFF,0xFF,0xFF,       //0x08
        0x00,0x00,0x00,0x00,0x00,0x3C,0x66,0x42,0x42,0x66,0x3C,0x00,0x00,0x00,0x00,0x00,       //0x09
        0xFF,0xFF,0xFF,0xFF,0xFF,0xC3,0x99,0xBD,0xBD,0x99,0xC3,0xFF,0xFF,0xFF,0xFF,0xFF,       //0x0A
        0x00,0x00,0x1E,0x0E,0x1A,0x32,0x78,0xCC,0xCC,0xCC,0xCC,0x78,0x00,0x00,0x00,0x00,       //0x0B
        0x00,0x00,0x3C,0x66,0x66,0x66,0x66,0x3C,0x18,0x7E,0x18,0x18,0x00,0x00,0x00,0x00,       //0x0C
        0x00,0x00,0x3F,0x33,0x3F,0x30,0x30,0x30,0x30,0x70,0xF0,0xE0,0x00,0x00,0x00,0x00,       //0x0D
        0x00,0x00,0x7F,0x63,0x7F,0x63,0x63,0x63,0x63,0x67,0xE7,0xE6,0xC0,0x00,0x00,0x00,       //0x0E
        0x00,0x00,0x00,0x18,0x18,0xDB,0x3C,0xE7,0x3C,0xDB,0x18,0x18,0x00,0x00,0x00,0x00,       //0x0F
        0x00,0x80,0xC0,0xE0,0xF0,0xF8,0xFE,0xF8,0xF0,0xE0,0xC0,0x80,0x00,0x00,0x00,0x00,       //0x10
        0x00,0x02,0x06,0x0E,0x1E,0x3E,0xFE,0x3E,0x1E,0x0E,0x06,0x02,0x00,0x00,0x00,0x00,       //0x11
        0x00,0x00,0x18,0x3C,0x7E,0x18,0x18,0x18,0x7E,0x3C,0x18,0x00,0x00,0x00,0x00,0x00,       //0x12
        0x00,0x00,0x66,0x66,0x66,0x66,0x66,0x66,0x66,0x00,0x66,0x66,0x00,0x00,0x00,0x00,       //0x13
        0x00,0x00,0x7F,0xDB,0xDB,0xDB,0x7B,0x1B,0x1B,0x1B,0x1B,0x1B,0x00,0x00,0x00,0x00,       //0x14
        0x00,0x7C,0xC6,0x60,0x38,0x6C,0xC6,0xC6,0x6C,0x38,0x0C,0xC6,0x7C,0x00,0x00,0x00,       //0x15
        0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0xFE,0xFE,0xFE,0xFE,0x00,0x00,0x00,0x00,       //0x16
        0x00,0x00,0x18,0x3C,0x7E,0x18,0x18,0x18,0x7E,0x3C,0x18,0x7E,0x00,0x00,0x00,0x00,       //0x17
        0x00,0x00,0x18,0x3C,0x7E,0x18,0x18,0x18,0x18,0x18,0x18,0x18,0x00,0x00,0x00,0x00,       //0x18
        0x00,0x00,0x18,0x18,0x18,0x18,0x18,0x18,0x18,0x7E,0x3C,0x18,0x00,0x00,0x00,0x00,       //0x19
        0x00,0x00,0x00,0x00,0x00,0x18,0x0C,0xFE,0x0C,0x18,0x00,0x00,0x00,0x00,0x00,0x00,       //0x1A
        0x00,0x00,0x00,0x00,0x00,0x30,0x60,0xFE,0x60,0x30,0x00,0x00,0x00,0x00,0x00,0x00,       //0x1B
        0x00,0x00,0x00,0x00,0x00,0x00,0xC0,0xC0,0xC0,0xFE,0x00,0x00,0x00,0x00,0x00,0x00,       //0x1C
        0x00,0x00,0x00,0x00,0x00,0x28,0x6C,0xFE,0x6C,0x28,0x00,0x00,0x00,0x00,0x00,0x00,       //0x1D
        0x00,0x00,0x00,0x00,0x10,0x38,0x38,0x7C,0x7C,0xFE,0xFE,0x00,0x00,0x00,0x00,0x00,       //0x1E
        0x00,0x00,0x00,0x00,0xFE,0xFE,0x7C,0x7C,0x38,0x38,0x10,0x00,0x00,0x00,0x00,0x00,       //0x1F
        0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,       //0x20' '
        0x00,0x00,0x18,0x3C,0x3C,0x3C,0x18,0x18,0x18,0x00,0x18,0x18,0x00,0x00,0x00,0x00,       //0x21'!'
        0x00,0x66,0x66,0x66,0x24,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,       //0x22'"'
        0x00,0x00,0x00,0x6C,0x6C,0xFE,0x6C,0x6C,0x6C,0xFE,0x6C,0x6C,0x00,0x00,0x00,0x00,       //0x23'#'
        0x18,0x18,0x7C,0xC6,0xC2,0xC0,0x7C,0x06,0x06,0x86,0xC6,0x7C,0x18,0x18,0x00,0x00,       //0x24'$'
        0x00,0x00,0x00,0x00,0xC2,0xC6,0x0C,0x18,0x30,0x60,0xC6,0x86,0x00,0x00,0x00,0x00,       //0x25'%'
        0x00,0x00,0x38,0x6C,0x6C,0x38,0x76,0xDC,0xCC,0xCC,0xCC,0x76,0x00,0x00,0x00,0x00,       //0x26'&'
        0x00,0x30,0x30,0x30,0x60,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,       //0x27'''
        0x00,0x00,0x0C,0x18,0x30,0x30,0x30,0x30,0x30,0x30,0x18,0x0C,0x00,0x00,0x00,0x00,       //0x28'('
        0x00,0x00,0x30,0x18,0x0C,0x0C,0x0C,0x0C,0x0C,0x0C,0x18,0x30,0x00,0x00,0x00,0x00,       //0x29')'
        0x00,0x00,0x00,0x00,0x00,0x66,0x3C,0xFF,0x3C,0x66,0x00,0x00,0x00,0x00,0x00,0x00,       //0x2A'*'
        0x00,0x00,0x00,0x00,0x00,0x18,0x18,0x7E,0x18,0x18,0x00,0x00,0x00,0x00,0x00,0x00,       //0x2B'+'
        0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x18,0x18,0x18,0x30,0x00,0x00,0x00,       //0x2C','
        0x00,0x00,0x00,0x00,0x00,0x00,0x00,0xFE,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,       //0x2D'-'
        0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x18,0x18,0x00,0x00,0x00,0x00,       //0x2E'.'
        0x00,0x00,0x00,0x00,0x02,0x06,0x0C,0x18,0x30,0x60,0xC0,0x80,0x00,0x00,0x00,0x00,       //0x2F'/'
        0x00,0x00,0x38,0x6C,0xC6,0xC6,0xD6,0xD6,0xC6,0xC6,0x6C,0x38,0x00,0x00,0x00,0x00,       //0x30'0'
        0x00,0x00,0x18,0x38,0x78,0x18,0x18,0x18,0x18,0x18,0x18,0x7E,0x00,0x00,0x00,0x00,       //0x31'1'
        0x00,0x00,0x7C,0xC6,0x06,0x0C,0x18,0x30,0x60,0xC0,0xC6,0xFE,0x00,0x00,0x00,0x00,       //0x32'2'
        0x00,0x00,0x7C,0xC6,0x06,0x06,0x3C,0x06,0x06,0x06,0xC6,0x7C,0x00,0x00,0x00,0x00,       //0x33'3'
        0x00,0x00,0x0C,0x1C,0x3C,0x6C,0xCC,0xFE,0x0C,0x0C,0x0C,0x1E,0x00,0x00,0x00,0x00,       //0x34'4'
        0x00,0x00,0xFE,0xC0,0xC0,0xC0,0xFC,0x06,0x06,0x06,0xC6,0x7C,0x00,0x00,0x00,0x00,       //0x35'5'
        0x00,0x00,0x38,0x60,0xC0,0xC0,0xFC,0xC6,0xC6,0xC6,0xC6,0x7C,0x00,0x00,0x00,0x00,       //0x36'6'
        0x00,0x00,0xFE,0xC6,0x06,0x06,0x0C,0x18,0x30,0x30,0x30,0x30,0x00,0x00,0x00,0x00,       //0x37'7'
        0x00,0x00,0x7C,0xC6,0xC6,0xC6,0x7C,0xC6,0xC6,0xC6,0xC6,0x7C,0x00,0x00,0x00,0x00,       //0x38'8'
        0x00,0x00,0x7C,0xC6,0xC6,0xC6,0x7E,0x06,0x06,0x06,0x0C,0x78,0x00,0x00,0x00,0x00,       //0x39'9'
        0x00,0x00,0x00,0x00,0x18,0x18,0x00,0x00,0x00,0x18,0x18,0x00,0x00,0x00,0x00,0x00,       //0x3A':'
        0x00,0x00,0x00,0x00,0x18,0x18,0x00,0x00,0x00,0x18,0x18,0x30,0x00,0x00,0x00,0x00,       //0x3B';'
        0x00,0x00,0x00,0x06,0x0C,0x18,0x30,0x60,0x30,0x18,0x0C,0x06,0x00,0x00,0x00,0x00,       //0x3C'<'
        0x00,0x00,0x00,0x00,0x00,0x7E,0x00,0x00,0x7E,0x00,0x00,0x00,0x00,0x00,0x00,0x00,       //0x3D'='
        0x00,0x00,0x00,0x60,0x30,0x18,0x0C,0x06,0x0C,0x18,0x30,0x60,0x00,0x00,0x00,0x00,       //0x3E'>'
        0x00,0x00,0x7C,0xC6,0xC6,0x0C,0x18,0x18,0x18,0x00,0x18,0x18,0x00,0x00,0x00,0x00,       //0x3F'?'
        0x00,0x00,0x00,0x7C,0xC6,0xC6,0xDE,0xDE,0xDE,0xDC,0xC0,0x7C,0x00,0x00,0x00,0x00,       //0x40'@'
        0x00,0x00,0x10,0x38,0x6C,0xC6,0xC6,0xFE,0xC6,0xC6,0xC6,0xC6,0x00,0x00,0x00,0x00,       //0x41'A'
        0x00,0x00,0xFC,0x66,0x66,0x66,0x7C,0x66,0x66,0x66,0x66,0xFC,0x00,0x00,0x00,0x00,       //0x42'B'
        0x00,0x00,0x3C,0x66,0xC2,0xC0,0xC0,0xC0,0xC0,0xC2,0x66,0x3C,0x00,0x00,0x00,0x00,       //0x43'C'
        0x00,0x00,0xF8,0x6C,0x66,0x66,0x66,0x66,0x66,0x66,0x6C,0xF8,0x00,0x00,0x00,0x00,       //0x44'D'
        0x00,0x00,0xFE,0x66,0x62,0x68,0x78,0x68,0x60,0x62,0x66,0xFE,0x00,0x00,0x00,0x00,       //0x45'E'
        0x00,0x00,0xFE,0x66,0x62,0x68,0x78,0x68,0x60,0x60,0x60,0xF0,0x00,0x00,0x00,0x00,       //0x46'F'
        0x00,0x00,0x3C,0x66,0xC2,0xC0,0xC0,0xDE,0xC6,0xC6,0x66,0x3A,0x00,0x00,0x00,0x00,       //0x47'G'
        0x00,0x00,0xC6,0xC6,0xC6,0xC6,0xFE,0xC6,0xC6,0xC6,0xC6,0xC6,0x00,0x00,0x00,0x00,       //0x48'H'
        0x00,0x00,0x3C,0x18,0x18,0x18,0x18,0x18,0x18,0x18,0x18,0x3C,0x00,0x00,0x00,0x00,       //0x49'I'
        0x00,0x00,0x1E,0x0C,0x0C,0x0C,0x0C,0x0C,0xCC,0xCC,0xCC,0x78,0x00,0x00,0x00,0x00,       //0x4A'J'
        0x00,0x00,0xE6,0x66,0x66,0x6C,0x78,0x78,0x6C,0x66,0x66,0xE6,0x00,0x00,0x00,0x00,       //0x4B'K'
        0x00,0x00,0xF0,0x60,0x60,0x60,0x60,0x60,0x60,0x62,0x66,0xFE,0x00,0x00,0x00,0x00,       //0x4C'L'
        0x00,0x00,0xC6,0xEE,0xFE,0xFE,0xD6,0xC6,0xC6,0xC6,0xC6,0xC6,0x00,0x00,0x00,0x00,       //0x4D'M'
        0x00,0x00,0xC6,0xE6,0xF6,0xFE,0xDE,0xCE,0xC6,0xC6,0xC6,0xC6,0x00,0x00,0x00,0x00,       //0x4E'N'
        0x00,0x00,0x7C,0xC6,0xC6,0xC6,0xC6,0xC6,0xC6,0xC6,0xC6,0x7C,0x00,0x00,0x00,0x00,       //0x4F'O'
        0x00,0x00,0xFC,0x66,0x66,0x66,0x7C,0x60,0x60,0x60,0x60,0xF0,0x00,0x00,0x00,0x00,       //0x50'P'
        0x00,0x00,0x7C,0xC6,0xC6,0xC6,0xC6,0xC6,0xC6,0xD6,0xDE,0x7C,0x0C,0x0E,0x00,0x00,       //0x51'Q'
        0x00,0x00,0xFC,0x66,0x66,0x66,0x7C,0x6C,0x66,0x66,0x66,0xE6,0x00,0x00,0x00,0x00,       //0x52'R'
        0x00,0x00,0x7C,0xC6,0xC6,0x60,0x38,0x0C,0x06,0xC6,0xC6,0x7C,0x00,0x00,0x00,0x00,       //0x53'S'
        0x00,0x00,0x7E,0x7E,0x5A,0x18,0x18,0x18,0x18,0x18,0x18,0x3C,0x00,0x00,0x00,0x00,       //0x54'T'
        0x00,0x00,0xC6,0xC6,0xC6,0xC6,0xC6,0xC6,0xC6,0xC6,0xC6,0x7C,0x00,0x00,0x00,0x00,       //0x55'U'
        0x00,0x00,0xC6,0xC6,0xC6,0xC6,0xC6,0xC6,0xC6,0x6C,0x38,0x10,0x00,0x00,0x00,0x00,       //0x56'V'
        0x00,0x00,0xC6,0xC6,0xC6,0xC6,0xD6,0xD6,0xD6,0xFE,0xEE,0x6C,0x00,0x00,0x00,0x00,       //0x57'W'
        0x00,0x00,0xC6,0xC6,0x6C,0x7C,0x38,0x38,0x7C,0x6C,0xC6,0xC6,0x00,0x00,0x00,0x00,       //0x58'X'
        0x00,0x00,0x66,0x66,0x66,0x66,0x3C,0x18,0x18,0x18,0x18,0x3C,0x00,0x00,0x00,0x00,       //0x59'Y'
        0x00,0x00,0xFE,0xC6,0x86,0x0C,0x18,0x30,0x60,0xC2,0xC6,0xFE,0x00,0x00,0x00,0x00,       //0x5A'Z'
        0x00,0x00,0x3C,0x30,0x30,0x30,0x30,0x30,0x30,0x30,0x30,0x3C,0x00,0x00,0x00,0x00,       //0x5B'['
        0x00,0x00,0x00,0x80,0xC0,0xE0,0x70,0x38,0x1C,0x0E,0x06,0x02,0x00,0x00,0x00,0x00,       //0x5C'\'
        0x00,0x00,0x3C,0x0C,0x0C,0x0C,0x0C,0x0C,0x0C,0x0C,0x0C,0x3C,0x00,0x00,0x00,0x00,       //0x5D']'
        0x10,0x38,0x6C,0xC6,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,       //0x5E'^'
        0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0xFF,0x00,0x00,       //0x5F'_'
        0x30,0x30,0x18,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,       //0x60'`'
        0x00,0x00,0x00,0x00,0x00,0x78,0x0C,0x7C,0xCC,0xCC,0xCC,0x76,0x00,0x00,0x00,0x00,       //0x61'a'
        0x00,0x00,0xE0,0x60,0x60,0x78,0x6C,0x66,0x66,0x66,0x66,0x7C,0x00,0x00,0x00,0x00,       //0x62'b'
        0x00,0x00,0x00,0x00,0x00,0x7C,0xC6,0xC0,0xC0,0xC0,0xC6,0x7C,0x00,0x00,0x00,0x00,       //0x63'c'
        0x00,0x00,0x1C,0x0C,0x0C,0x3C,0x6C,0xCC,0xCC,0xCC,0xCC,0x76,0x00,0x00,0x00,0x00,       //0x64'd'
        0x00,0x00,0x00,0x00,0x00,0x7C,0xC6,0xFE,0xC0,0xC0,0xC6,0x7C,0x00,0x00,0x00,0x00,       //0x65'e'
        0x00,0x00,0x38,0x6C,0x64,0x60,0xF0,0x60,0x60,0x60,0x60,0xF0,0x00,0x00,0x00,0x00,       //0x66'f'
        0x00,0x00,0x00,0x00,0x00,0x76,0xCC,0xCC,0xCC,0xCC,0xCC,0x7C,0x0C,0xCC,0x78,0x00,       //0x67'g'
        0x00,0x00,0xE0,0x60,0x60,0x6C,0x76,0x66,0x66,0x66,0x66,0xE6,0x00,0x00,0x00,0x00,       //0x68'h'
        0x00,0x00,0x18,0x18,0x00,0x38,0x18,0x18,0x18,0x18,0x18,0x3C,0x00,0x00,0x00,0x00,       //0x69'i'
        0x00,0x00,0x06,0x06,0x00,0x0E,0x06,0x06,0x06,0x06,0x06,0x06,0x66,0x66,0x3C,0x00,       //0x6A'j'
        0x00,0x00,0xE0,0x60,0x60,0x66,0x6C,0x78,0x78,0x6C,0x66,0xE6,0x00,0x00,0x00,0x00,       //0x6B'k'
        0x00,0x00,0x38,0x18,0x18,0x18,0x18,0x18,0x18,0x18,0x18,0x3C,0x00,0x00,0x00,0x00,       //0x6C'l'
        0x00,0x00,0x00,0x00,0x00,0xEC,0xFE,0xD6,0xD6,0xD6,0xD6,0xC6,0x00,0x00,0x00,0x00,       //0x6D'm'
        0x00,0x00,0x00,0x00,0x00,0xDC,0x66,0x66,0x66,0x66,0x66,0x66,0x00,0x00,0x00,0x00,       //0x6E'n'
        0x00,0x00,0x00,0x00,0x00,0x7C,0xC6,0xC6,0xC6,0xC6,0xC6,0x7C,0x00,0x00,0x00,0x00,       //0x6F'o'
        0x00,0x00,0x00,0x00,0x00,0xDC,0x66,0x66,0x66,0x66,0x66,0x7C,0x60,0x60,0xF0,0x00,       //0x70'p'
        0x00,0x00,0x00,0x00,0x00,0x76,0xCC,0xCC,0xCC,0xCC,0xCC,0x7C,0x0C,0x0C,0x1E,0x00,       //0x71'q'
        0x00,0x00,0x00,0x00,0x00,0xDC,0x76,0x66,0x60,0x60,0x60,0xF0,0x00,0x00,0x00,0x00,       //0x72'r'
        0x00,0x00,0x00,0x00,0x00,0x7C,0xC6,0x60,0x38,0x0C,0xC6,0x7C,0x00,0x00,0x00,0x00,       //0x73's'
        0x00,0x00,0x10,0x30,0x30,0xFC,0x30,0x30,0x30,0x30,0x36,0x1C,0x00,0x00,0x00,0x00,       //0x74't'
        0x00,0x00,0x00,0x00,0x00,0xCC,0xCC,0xCC,0xCC,0xCC,0xCC,0x76,0x00,0x00,0x00,0x00,       //0x75'u'
        0x00,0x00,0x00,0x00,0x00,0x66,0x66,0x66,0x66,0x66,0x3C,0x18,0x00,0x00,0x00,0x00,       //0x76'v'
        0x00,0x00,0x00,0x00,0x00,0xC6,0xC6,0xD6,0xD6,0xD6,0xFE,0x6C,0x00,0x00,0x00,0x00,       //0x77'w'
        0x00,0x00,0x00,0x00,0x00,0xC6,0x6C,0x38,0x38,0x38,0x6C,0xC6,0x00,0x00,0x00,0x00,       //0x78'x'
        0x00,0x00,0x00,0x00,0x00,0xC6,0xC6,0xC6,0xC6,0xC6,0xC6,0x7E,0x06,0x0C,0xF8,0x00,       //0x79'y'
        0x00,0x00,0x00,0x00,0x00,0xFE,0xCC,0x18,0x30,0x60,0xC6,0xFE,0x00,0x00,0x00,0x00,       //0x7A'z'
        0x00,0x00,0x0E,0x18,0x18,0x18,0x70,0x18,0x18,0x18,0x18,0x0E,0x00,0x00,0x00,0x00,       //0x7B'{'
        0x00,0x00,0x18,0x18,0x18,0x18,0x00,0x18,0x18,0x18,0x18,0x18,0x00,0x00,0x00,0x00,       //0x7C'|'
        0x00,0x00,0x70,0x18,0x18,0x18,0x0E,0x18,0x18,0x18,0x18,0x70,0x00,0x00,0x00,0x00,       //0x7D'}'
        0x00,0x00,0x76,0xDC,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,       //0x7E'~'
        0x00,0x00,0x00,0x00,0x10,0x38,0x6C,0xC6,0xC6,0xC6,0xFE,0x00,0x00,0x00,0x00,0x00,       //0x7F''
        0x00,0x00,0x3C,0x66,0xC2,0xC0,0xC0,0xC0,0xC2,0x66,0x3C,0x0C,0x06,0x7C,0x00,0x00,       //0x80
        0x00,0x00,0xCC,0x00,0x00,0xCC,0xCC,0xCC,0xCC,0xCC,0xCC,0x76,0x00,0x00,0x00,0x00,       //0x81
        0x00,0x0C,0x18,0x30,0x00,0x7C,0xC6,0xFE,0xC0,0xC0,0xC6,0x7C,0x00,0x00,0x00,0x00,       //0x82
        0x00,0x10,0x38,0x6C,0x00,0x78,0x0C,0x7C,0xCC,0xCC,0xCC,0x76,0x00,0x00,0x00,0x00,       //0x83
        0x00,0x00,0xCC,0x00,0x00,0x78,0x0C,0x7C,0xCC,0xCC,0xCC,0x76,0x00,0x00,0x00,0x00,       
    };


    //////////////////////////////////////////////////////////////////
    // 功能： 产生 25MHz 的像素时钟 R_clk_25M
    //////////////////////////////////////////////////////////////////
    always @(posedge I_clk or negedge I_rst_n) // 输入的 50 MHz I_clk 的上升沿
    begin
        if(!I_rst_n) // reset
            R_clk_25M   <=  1'b0        ;
        else
            R_clk_25M   <=  ~R_clk_25M  ;     // 每到上升沿才反转，50 MHz -> 25 MHz
    end

    //////////////////////////////////////////////////////////////////
    // 功能：产生行时序计数器 R_h_cnt
    //////////////////////////////////////////////////////////////////
    always @(posedge R_clk_25M or negedge I_rst_n)
    begin
        if(!I_rst_n) // reset
            R_h_cnt <=  12'd0   ;
        else if(R_h_cnt == C_H_LINE_PERIOD - 1'b1) // 计数到最大值了，重新开始
            R_h_cnt <=  12'd0   ;
        else
            R_h_cnt <=  R_h_cnt + 1'b1  ;                
    end                

    // 产生行时序输出 O_hs，C_H_SYNC_PULSE 内要置零
    assign O_hs =   (R_h_cnt < C_H_SYNC_PULSE) ? 1'b0 : 1'b1    ; 
    //////////////////////////////////////////////////////////////////


    //////////////////////////////////////////////////////////////////
    // 功能：产生场时序计数器 R_v_cnt
    //////////////////////////////////////////////////////////////////
    always @(posedge R_clk_25M or negedge I_rst_n)
    begin
        if(!I_rst_n) // reset
            R_v_cnt <=  12'd0   ;
        else if(R_v_cnt == C_V_FRAME_PERIOD - 1'b1) // 计数到最大值了，重新开始
            R_v_cnt <=  12'd0   ;
        else if(R_h_cnt == C_H_LINE_PERIOD - 1'b1) // 一行完成了，R_v_cnt++
            R_v_cnt <=  R_v_cnt + 1'b1  ;
        else // 不变
            R_v_cnt <=  R_v_cnt ;                        
    end                

    // 产生行时序输出 O_vs，C_V_SYNC_PULSE 内要置零
    assign O_vs =   (R_v_cnt < C_V_SYNC_PULSE) ? 1'b0 : 1'b1    ; 
    //////////////////////////////////////////////////////////////////  


    // 产生 是否可以输出 RGB: W_active_flag 
    // 可以输出：R_h_cnt 在行消隐、行前肩之间，且 R_v_cnt 在场消隐、场前肩之间
    assign W_active_flag =  (R_h_cnt >= (C_H_SYNC_PULSE + C_H_BACK_PORCH                  ))  &&
                            (R_h_cnt <= (C_H_SYNC_PULSE + C_H_BACK_PORCH + C_H_ACTIVE_TIME))  && 
                            (R_v_cnt >= (C_V_SYNC_PULSE + C_V_BACK_PORCH                  ))  &&
                            (R_v_cnt <= (C_V_SYNC_PULSE + C_V_BACK_PORCH + C_V_ACTIVE_TIME))  ;  
    //////////////////////////////////////////////////////////////////                     


    //////////////////////////////////////////////////////////////////
    // 功能：在 VGA 显示屏上同步 shell 的输出内容
    //////////////////////////////////////////////////////////////////
    always @(posedge R_clk_25M or negedge I_rst_n)
    begin
        if(!I_rst_n) // reset
            begin
                O_red   <=  4'b0000   ;
                O_green <=  4'b0000   ;
                O_blue  <=  4'b0000   ; 
            end
        else if(W_active_flag)     // 如果现在可以输出 RGB
            begin
                // 得到当前字符的 x 坐标
                R_char_h_cnt    <=  (R_h_cnt - C_H_SYNC_PULSE - C_H_BACK_PORCH) / 10 ;
                // 得到当前字符的 y 坐标
                R_char_v_cnt    <=  (R_v_cnt - C_V_SYNC_PULSE - C_V_BACK_PORCH) / 20 ;
                // 得到当前字符的 8 位 ascii 码
                R_now_ascii     <=  I_string[8 * (R_char_v_cnt * 64 + R_char_h_cnt + 1) - : 8]  ;
                // 得到当前字符 字模的 x 坐标
                R_char_h_detail <=  R_h_cnt - C_H_SYNC_PULSE - C_H_BACK_PORCH - R_char_h_cnt * 10;
                // 得到当前字符 字模的 y 坐标
                R_char_v_detail <=  R_v_cnt - C_V_SYNC_PULSE - C_V_BACK_PORCH - R_char_v_cnt * 20;

                // 取字模
                if(R_char_h_detail < 1 || R_char_h_detail >= 9 || R_char_v_detail < 2 || R_char_v_detail >= 18)
                    begin // 因为我们的像素是 10 * 20，而字模是 8 * 16，所以边缘不输出
                        O_red   <=  4'b0000   ;
                        O_green <=  4'b0000   ;
                        O_blue  <=  4'b0000   ; 
                    end  
                else if(C_ascii_character[R_now_ascii * 16 + R_char_v_detail - 2][R_char_h_detail - 1] == 1)
                    begin // 要输出的，全白，全 1
                        O_red   <=  4'b1111    ;
                        O_green <=  4'b1111    ;
                        O_blue  <=  4'b1111    ;
                    end
                else
                    begin
                        O_red   <=  4'b0000   ;
                        O_green <=  4'b0000   ;
                        O_blue  <=  4'b0000   ; 
                    end  
            end
        else // 现在不能输出 RGB
            begin
                O_red   <=  4'b0000    ;
                O_green <=  4'b0000    ;
                O_blue  <=  4'b0000    ; 
            end           
    end

        
endmodule




